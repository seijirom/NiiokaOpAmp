* Z:\HOME\ANAGIX\WORK\2020SEPTO\NIIOKAOPAMP\OAMP_KLAYOUT_TB.ASC
*V1 N001 0 5
*XX1 N003 N002 N001 N001 N002 0 OPAMP_K_NIIOKA_20200903
*V2 N003 0 2.5 AC 1 0
*
* BLOCK SYMBOL DEFINITIONS
.SUBCKT OPAMP_K_NIIOKA_20200903 IN+ IN_ VB VDD OUT GND
M1 N002 N001 VDD VDD PMOS L=3U W=100U
M2 N001 N001 VDD VDD PMOS L=3U W=100U
M4 N001 IN_ N004 GND NMOS L=1U W=400U
M5 N002 IN+ N004 GND NMOS L=1U W=400U
M6 N004 N003 GND GND NMOS L=2.5U W=120U
M7 N003 N003 GND GND NMOS L=2.5U W=10U
M8 OUT N003 GND GND NMOS L=1U W=120U
M3 OUT N002 VDD VDD PMOS L=1U W=240U
R1 N003 VB 40K
C2 N002 N001 3P
*.INCLUDE "./MODELS/OR1_MOS"
.ENDS OPAMP_K_NIIOKA_20200903

.MODEL NMOS NMOS
.MODEL PMOS PMOS
.LIB C:\USERS\ANAGIX\MY DOCUMENTS\LTSPICEXVII\LIB\CMP\STANDARD.MOS
*.INCLUDE "./MODELS/OR1_MOS"
.AC DEC 100 1 1G
.BACKANNO
.END
