* Z:\HOME\ANAGIX\WORK\2020SEPTO\NIIOKAOPAMP\OPAMP_K_NIIOKA_20200903.ASC
M1 N002 N001 VDD VDD PCH L=3U W=100U
M2 N001 N001 VDD VDD PCH L=3U W=100U
M4 N001 IN+ N004 0 NCH L=1U W=400U
M5 N002 IN_ N004 0 NCH L=1U W=400U
M6 N004 N003 0 0 NCH L=2.5U W=120U
M7 N003 N003 0 0 NCH L=2.5U W=10U
M8 OUT N003 0 0 NCH L=1U W=120U
M3 OUT N002 VDD VDD PCH L=1U W=240U
C1 N002 OUT 3.0264P
R1 N003 VB 4K
.MODEL NMOS NMOS
.MODEL PMOS PMOS
.LIB C:\USERS\ANAGIX\MY DOCUMENTS\LTSPICEXVII\LIB\CMP\STANDARD.MOS
*.INCLUDE "./MODELS/OR1_MOS"
.TRAN 10M
.BACKANNO
.END
