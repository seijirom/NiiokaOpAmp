* Created by KLayout

* cell niioka_new
.SUBCKT niioka_new
* net 1 Vb
* net 2 Vdd
* net 4 Vout
* net 8 Vin+
* net 9 Vin-
* net 10 Vss
* device instance $1 r0 *1 198,319.75 CAP
C$1 5 6 3.0264e-12
* device instance $2 r0 *1 65.5,322 HRES
R$2 3 1 40250
* device instance $3 r0 *1 49.75,293 NMOS
M$3 10 3 3 10 NMOS L=2.5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $4 r180 *1 166.5,315.5 PMOS
M$4 4 6 2 2 PMOS L=1U W=240U AS=280P AD=280P PS=294U PD=294U
* device instance $10 r0 *1 154,269.5 NMOS
M$10 10 3 4 10 NMOS L=1U W=120U AS=144P AD=144P PS=156U PD=156U
* device instance $15 r180 *1 93.5,323.5 PMOS
M$15 5 5 2 2 PMOS L=3U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $19 m0 *1 115,323.5 PMOS
M$19 6 5 2 2 PMOS L=3U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $23 r180 *1 96,277 NMOS
M$23 5 8 7 10 NMOS L=1U W=400U AS=440P AD=440P PS=462U PD=462U
* device instance $33 r180 *1 136.5,277 NMOS
M$33 6 9 7 10 NMOS L=1U W=400U AS=440P AD=440P PS=462U PD=462U
* device instance $43 r180 *1 54.75,267 NMOS
M$43 7 3 10 10 NMOS L=2.5U W=120U AS=140P AD=140P PS=154U PD=154U
.ENDS niioka_new
